package NocConstants is
end package;